parameter DWIDTH  = 16;
parameter INSIZE  = 12;
parameter FSIZE   = 5;
parameter PSIZE   = 2;
parameter N_F1    = 20;
parameter N_F2    = 50;
parameter OUTSIZE = 10;
parameter WSIZE   = 13;
parameter IFMSIZE = 9;
parameter FACCUM  = 7;
parameter PACCUM  = 8;
parameter LWIDTH  = 8;
parameter STEP    = 10;
