../src/parameters.vh